module alu (input [7:0] regA, regB,
				input [1:0] opcode,
				input clock, computestrobe,
				output reg [7:0] result;
				);

				
	always @(posedge clock) begin
		if (computestrobe) begin 
			
			
			
			
			
		end
	end


endmodule 