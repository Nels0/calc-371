module calculator ()



endmodule 